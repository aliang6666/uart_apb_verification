package apb_agent_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "param_def.v"


`include "reg_trans.sv"
`include "reg_driver.sv"
`include "reg_monitor.sv"
`include "reg_sequence.sv"
`include "reg_sequencer.sv"
`include "reg_agent.sv"
endpackage